----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 27.01.2016 23:26:13
-- Design Name: 
-- Module Name: KSAred - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity KSAred is
    Port ( A : in STD_LOGIC;
           B : in STD_LOGIC;
           P : out STD_LOGIC;
           G : out STD_LOGIC);
end KSAred;

architecture Behavioral of KSAred is
begin

    P <= A xor B;
    G <= A and B;

end Behavioral;
